library verilog;
use verilog.vl_types.all;
entity clk is
    port(
        c7              : out    vl_logic;
        pin_name1       : in     vl_logic;
        a1              : out    vl_logic;
        b1              : out    vl_logic;
        d1              : out    vl_logic;
        e1              : out    vl_logic;
        f1              : out    vl_logic;
        g1              : out    vl_logic;
        a0              : out    vl_logic;
        b0              : out    vl_logic;
        c0              : out    vl_logic;
        d0              : out    vl_logic;
        e0              : out    vl_logic;
        f0              : out    vl_logic;
        g0              : out    vl_logic;
        a               : out    vl_logic;
        b               : out    vl_logic;
        c               : out    vl_logic;
        d               : out    vl_logic;
        e               : out    vl_logic;
        f               : out    vl_logic;
        g               : out    vl_logic
    );
end clk;
