library verilog;
use verilog.vl_types.all;
entity clk_vlg_check_tst is
    port(
        a               : in     vl_logic;
        a0              : in     vl_logic;
        a1              : in     vl_logic;
        b               : in     vl_logic;
        b0              : in     vl_logic;
        b1              : in     vl_logic;
        c               : in     vl_logic;
        c0              : in     vl_logic;
        c7              : in     vl_logic;
        d               : in     vl_logic;
        d0              : in     vl_logic;
        d1              : in     vl_logic;
        e               : in     vl_logic;
        e0              : in     vl_logic;
        e1              : in     vl_logic;
        f               : in     vl_logic;
        f0              : in     vl_logic;
        f1              : in     vl_logic;
        g               : in     vl_logic;
        g0              : in     vl_logic;
        g1              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end clk_vlg_check_tst;
