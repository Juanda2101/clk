library verilog;
use verilog.vl_types.all;
entity clk_vlg_sample_tst is
    port(
        pin_name1       : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end clk_vlg_sample_tst;
